// https://hdlbits.01xz.net/wiki/Exams/2012_q1g

module top_module (
    input [4:1] x,
    output f );

    // sum of product
    // assign f = (~x[2] & ~x[4]) | (~x[1] & x[3]) | (x[2] & x[3] & x[4]);

    // product of sum
    assign f = (x[3] | ~x[4]) & (~x[2] | x[3]) & (~x[1] | ~x[2] | x[4]) & (~x[1] | x[2] | ~x[4]);

endmodule

