// https://hdlbits.01xz.net/wiki/Exams/m2014_q4h

module top_module (
    input in,
    output out);

    assign out = in;
endmodule
