/***********************************************************************************************
FILE NAME           module1.v
DEPARTMENT          Logic
AUTHOR              XU Lu
AUTHOR'S EMAIL      xu.lu@tnc.ltd
------------------------------------------------------------------------------------------------
RELEASE HISTORY
VERSION             DATE            AUTHOR      DESCRIPTION
1.0                 2024-06-28      XU Lu       Initial
------------------------------------------------------------------------------------------------
KEYWORDS            pre process, sync word
------------------------------------------------------------------------------------------------
PURPOSE             use for match sync word and output frame data with defined length
***********************************************************************************************/

/**********************************************************************************************
MODULE DEFINITION
**********************************************************************************************/
`timescale  1ns / 1ps
module module1 (
    // RESET & CLOCK
    input  wire clk,
    input  wire rstn,
    // IN INTERFACE
    input  wire in,
    // OUTPUT INTERFACE
    output reg out
);

    /***************************************
        PARAMETER SEGMENT
    ***************************************/

    /***************************************
        WIRE SEGMENT
    ***************************************/

    /***************************************
        REGISTER SEGMENT
    ***************************************/

    /***************************************
        INSTANCE SEGMENT
    ***************************************/

    /***************************************
        ASSIGN SEGMENT
    ***************************************/

    /***************************************
        ALWAYS SEGMENT
    ***************************************/
    always @(posedge clk) begin
        if(~rstn) begin
            out <= 1'b0;
        end else begin
            out <= in;
        end
    end

endmodule // <--- module1 module end
