// https://hdlbits.01xz.net/wiki/Exams/m2014_q4i

module top_module (
    output out);

    assign out = 1'b0;
endmodule
